module Tester;

integer i;
real k;

initial
begin
	for (i = 0; 1 === 1; i++)
	begin
		k = k * k;
		$display("tester");
	end

	$finish;
end


initial
begin
	for (i = 0; 1 === 1; i++)
	begin
		k = k * k;
		$display("tester");
	end

	$finish;
end


initial
begin
	for (i = 0; 1 === 1; i++)
	begin
		k = k * k;
		$display("tester");
	end

	$finish;
end


initial
begin
	for (i = 0; 1 === 1; i++)
	begin
		k = k * k;
		$display("tester");
	end

	$finish;
end
endmodule
